package fifo_pkg;
  import uvm_pkg::*;
`include "uvm_macros.svh"
// `include "test.sv"
`include "fifo_parameter.sv"
`include "fifo_seq_item.sv"
`include "fifo_sequence.sv"
`include "fifo_sequencer.sv"
`include "fifo_driver.sv"
`include "fifo_imon.sv"
`include "fifo_omon.sv"
`include "fifo_scoreboard.sv"
`include "master_agent.sv"
`include "slave_agent.sv"
`include "fifo_env.sv"
// `include "fifo_subscriber.sv"

endpackage
  
