typedef uvm_sequencer#(transaction) sequencer;