parameter DATA_WIDTH=8;
parameter ADDR_WIDTH=5;
parameter ADDR_BUS_WIDTH=4; 	
parameter MEM_SIZE=31;
